module ImageGenerator (readyToBeProcessed, encryptedSubmatrixElements, processed);
input readyToBeProcessed;
input [15:0] encryptedSubmatrixElements;
output processed;

endmodule

