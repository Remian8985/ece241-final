module ece241final();


endmodule 