//Uses the AES encryption algorithm to encrypt 160 by 120 pixel
//Displays the encrypted image via VGA
module ImageEncryptor;

endmodule 

